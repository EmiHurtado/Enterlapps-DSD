library ieee;
use ieee.std_logic_1164.all;

entity ConvertidorVectorUnitario8 is
	port(
		a, b, c, d, e, f, g, h : out std_logic;
		entradaVector : in std_logic_vector(0 to 7)
	);
end ConvertidorVectorUnitario8; 

architecture ConvVecUni8 of ConvertidorVectorUnitario8 is

begin
	a <= entradaVector(0);
	b <= entradaVector(1);
	c <= entradaVector(2);
	d <= entradaVector(3);
	e <= entradaVector(4);
	f <= entradaVector(5);
	g <= entradaVector(6);
	h <= entradaVector(7);
	
end ConvVecUni8;