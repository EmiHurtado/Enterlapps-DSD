library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity GeneradorVideo is
    port (
        CLK : in std_logic;
        
    );
end entity GeneradorVideo;