library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity RegCorrimiento3 is
	port (
	   CLK, RESET, CARGA : in std_logic;
		ENTRADA		: in std_logic_vector(7 downto 0);
		SALIDA		: out std_logic_vector(7 downto 0)
	);
end RegCorrimiento3;  

architecture funcion3 of RegCorrimiento3 is 
	signal REGISTRO 	: std_logic_vector(7 downto 0);
	signal contador	: integer range 0 to 8 := 0;

begin	 
	Multiplexor: process(CLK, RESET, CARGA, ENTRADA)
	begin
		--REGISTRO DE CORRIMIENTO: ENTRADA PARALELO/SALIDA SERIE, DESPLAZAMIENTO A LA DERECHA
	
							if RESET = '0' then
										REGISTRO <= (others => '0');
			
							elsif(CLK'event and CLK = '1') then
									if(CARGA = '1') then
										REGISTRO <= ENTRADA;
									else
										if(contador = 8) then
										contador <= 0;
										else
											REGISTRO(6 downto 0) <= REGISTRO(7 downto 1);
											contador <= contador + 1 ;
										end if;
									end if;
									
							end if;
		
	end process;
		SALIDA(0) <= REGISTRO(0);

end funcion3;